module bi_constants_rom (
    input [3:0] index,
    output reg signed [0:319] bi_yplus_x,
    output reg signed [0:319] bi_yminus_x,
    output reg signed [0:319] bi_z
);

    // ROM implementation using case statement
    always @(*) begin
        case(index)
            3'd0: begin
                bi_yplus_x = {
     32'd2047605, -32'd6079156, -32'd11754271, 32'd27544626, 32'd4014787, 
    -32'd12694345, 32'd3660896, 32'd29566456, -32'd14356035, 32'd25967493
    // Complete with zeros to make 320 bits
};
                bi_yminus_x = {
    -32'd15469378, 32'd19500929, 32'd5043384, 32'd12720692, 32'd9406986, 
    -32'd727428, 32'd3049990, -32'd2722910, 32'd934262, -32'd12545711
    // Complete with zeros to make 320 bits
};

                bi_z = {
     -32'd4438546, -32'd24514362, 32'd11864899, 32'd29287919, -32'd12363380, 
    32'd10184609, -32'd14785194, 32'd9688441, 32'd4489570, -32'd8738181
    // Complete with zeros to make 320 bits
};
       end
            
            3'd1: begin
                bi_yplus_x = {
    -32'd1550024, 32'd28944400, -32'd14772189, 32'd27787600, -32'd16685262, 
    32'd616977, -32'd7912398, 32'd24204773, -32'd9688557, 32'd15636291
    // Complete with zeros to make 320 bits
};
                bi_yminus_x = {
    32'd11199574, 32'd7689662, -32'd11775962, 32'd16354577, -32'd11807043, 
    32'd15682896, -32'd1102322, -32'd11556148, 32'd4717097, 32'd16568933
    // Complete with zeros to make 320 bits
};
                bi_z = {
    -32'd9920357, -32'd17749093, 32'd10017326, 32'd7512774, 32'd15915852, 
    32'd23220365, -32'd15670865, -32'd11779434, -32'd5976125, 32'd30464156
    // Complete with zeros to make 320 bits
};
            end
            
            3'd2: begin
                bi_yplus_x = {
    32'd10819380, -32'd15438304, 32'd14515107, 32'd32867885, 32'd12577861, 
    -32'd30064349, 32'd1981175, 32'd27284546, 32'd11473154, 32'd10861363
    // Complete with zeros to make 320 bits
};
                bi_yminus_x = {
    32'd5581306, -32'd12668491, 32'd12483688, -32'd25653668, 32'd6594696, 
    -32'd11272109, 32'd9066809, 32'd20377586, 32'd6336745, 32'd4708026
    // Complete with zeros to make 320 bits
};
                bi_z = {
    -32'd15815942, -32'd23678021, 32'd13850243, 32'd28542350, -32'd4348115, 
    32'd10237984, 32'd4097519, -32'd29386857, 32'd16186464, 32'd19563160
    // Complete with zeros to make 320 bits
};
            end
            
            3'd3: begin
                bi_yplus_x = {
    -32'd15175766, -32'd23952439, 32'd5230134, 32'd19480852, 32'd5516873, 
    32'd30523605, -32'd2777874, 32'd1723747, 32'd9909285, 32'd5153746
    // Complete with zeros to make 320 bits
};
                bi_yminus_x = {
    32'd7715701, 32'd30598449, 32'd16520125, 32'd20654025, 32'd1649722, 
    32'd28475525, 32'd10083793, 32'd7665486, -32'd3463509, -32'd30269007
    // Complete with zeros to make 320 bits
};
                bi_z = {
    -32'd1409300, 32'd29794553, 32'd1370708, -32'd31400660, 32'd7843316, 
    -32'd20181635, 32'd3680757, 32'd9657904, 32'd14381568, 32'd28881845
    // Complete with zeros to make 320 bits
};
            end
            
            3'd4: begin
                bi_yplus_x = {
    32'd13821877, -32'd13062696, -32'd1361450, 32'd18474211, 32'd8844726, 
    -32'd23510406, -32'd8745502, 32'd14201702, -32'd6692182, -32'd22518993
    // Complete with zeros to make 320 bits
};
                bi_yminus_x = {
    -32'd14220951, 32'd18853322, -32'd7212327, 32'd31655028, -32'd10571707, 
    -32'd27098617, -32'd4740862, 32'd3374702, -32'd7839871, -32'd6455177
    // Complete with zeros to make 320 bits
};
                bi_z = {
    -32'd3209784, 32'd2207753, -32'd10431137, -32'd8514358, -32'd2830569, 
    -32'd7602672, -32'd12240689, -32'd28974889, -32'd12963868, 32'd4566830
    // Complete with zeros to make 320 bits
};
            end
            
            3'd5: begin
                bi_yplus_x = {
    -32'd16132436, -32'd31111463, -32'd663000, -32'd12437364, -32'd9423865, 
    -32'd6854661, 32'd7868801, 32'd29681144, -32'd4185821, -32'd25154831
    // Complete with zeros to make 320 bits
};
                bi_yminus_x = {
    32'd6466918, 32'd171356, 32'd15725684, 32'd3844789, 32'd9300885, 
    32'd16472782, -32'd11814844, 32'd7349804, -32'd2703214, 32'd25576264
    // Complete with zeros to make 320 bits
};
                bi_z = {
    32'd16193877, -32'd30714912, -32'd14088058, 32'd8965339, -32'd15038942, 
    32'd817875, -32'd16149481, 32'd9739013, 32'd13316479, 32'd23103977
    // Complete with zeros to make 320 bits
};
            end
            
            3'd6: begin
                bi_yplus_x = {
    32'd9256800, -32'd18074513, 32'd4729455, 32'd17238398, -32'd16270840, 
    -32'd16903474, 32'd14003687, -32'd2394130, 32'd3180713, -32'd33521811
    // Complete with zeros to make 320 bits
};
                bi_yminus_x = {
    32'd630305, -32'd19827198, 32'd9761698, 32'd22616405, 32'd11360617, 
    -32'd21236817, 32'd5036987, 32'd32336398, -32'd4174131, -32'd25182317
    // Complete with zeros to make 320 bits
};
                bi_z = {
    -32'd14291300, -32'd2449256, -32'd15960994, -32'd6554551, -32'd5774029, 
    32'd9494427, -32'd7406481, -32'd24237460, 32'd2639453, -32'd13720693
    // Complete with zeros to make 320 bits
};
            end
            
            3'd7: begin
                bi_yplus_x = {
    -32'd7894876, 32'd25105118, 32'd15033784, -32'd18940575, -32'd863023, 
    -32'd31907062, 32'd6866145, 32'd9282714, -32'd5046075, -32'd3151181
    // Complete with zeros to make 320 bits
};
                bi_yminus_x = {
    -32'd15804619, 32'd2198790, -32'd2625887, 32'd1573892, -32'd5090925, 
    -32'd11662737, -32'd14592823, -32'd31801215, 32'd15950226, -32'd24326370
    // Complete with zeros to make 320 bits
};
                bi_z = {
    -32'd12290683, -32'd32461234, -32'd16236442, -32'd13812022, -32'd2735503, 
    -32'd5446979, 32'd7453183, -32'd2241613, 32'd10324967, -32'd3099351
    // Complete with zeros to make 320 bits
};
            end
            
            default: begin
                bi_yplus_x = {320{1'b0}};
                bi_yminus_x = {320{1'b0}};
                bi_z = {320{1'b0}};
            end
        endcase
    end

endmodule
